`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/12/2023 12:48:57 AM
// Design Name: 
// Module Name: cybercobra
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CYBERcobra
(
    input  logic            clk_i,
    input  logic            rst_i,
    input  logic    [15:0]  sw_i,
    output logic    [31:0]  out_o
);
    
    

endmodule
